module led_rgb_pwm(
);

endmodule